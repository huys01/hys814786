
//----------------------------------------------------------------------------
// File : sine_lut64_14bit.vh
//----------------------------------------------------------------------------
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 
//
//----------------------------------------------------------------------------

  assign sine_lut64_14bit[0]  = 14'h2000;
  assign sine_lut64_14bit[1]  = 14'h2322;
  assign sine_lut64_14bit[2]  = 14'h263D;
  assign sine_lut64_14bit[3]  = 14'h2949;
  assign sine_lut64_14bit[4]  = 14'h2C3E;
  assign sine_lut64_14bit[5]  = 14'h2F15;
  assign sine_lut64_14bit[6]  = 14'h31C6;
  assign sine_lut64_14bit[7]  = 14'h344C;
  assign sine_lut64_14bit[8]  = 14'h369F;
  assign sine_lut64_14bit[9]  = 14'h38BB;
  assign sine_lut64_14bit[10] = 14'h3A9A;
  assign sine_lut64_14bit[11] = 14'h3C37;
  assign sine_lut64_14bit[12] = 14'h3D8F;
  assign sine_lut64_14bit[13] = 14'h3E9E;
  assign sine_lut64_14bit[14] = 14'h3F61;
  assign sine_lut64_14bit[15] = 14'h3FD7;
  assign sine_lut64_14bit[16] = 14'h3FFF;
  assign sine_lut64_14bit[17] = 14'h3FD7;
  assign sine_lut64_14bit[18] = 14'h3F61;
  assign sine_lut64_14bit[19] = 14'h3E9E;
  assign sine_lut64_14bit[20] = 14'h3D8F;
  assign sine_lut64_14bit[21] = 14'h3C37;
  assign sine_lut64_14bit[22] = 14'h3A9A;
  assign sine_lut64_14bit[23] = 14'h38BB;
  assign sine_lut64_14bit[24] = 14'h369F;
  assign sine_lut64_14bit[25] = 14'h344C;
  assign sine_lut64_14bit[26] = 14'h31C6;
  assign sine_lut64_14bit[27] = 14'h2F15;
  assign sine_lut64_14bit[28] = 14'h2C3E;
  assign sine_lut64_14bit[29] = 14'h2949;
  assign sine_lut64_14bit[30] = 14'h263D;
  assign sine_lut64_14bit[31] = 14'h2322;
  assign sine_lut64_14bit[32] = 14'h2000;
  assign sine_lut64_14bit[33] = 14'h1CDD;
  assign sine_lut64_14bit[34] = 14'h19C2;
  assign sine_lut64_14bit[35] = 14'h16B6;
  assign sine_lut64_14bit[36] = 14'h13C1;
  assign sine_lut64_14bit[37] = 14'h10EA;
  assign sine_lut64_14bit[38] = 14'hE39;
  assign sine_lut64_14bit[39] = 14'hBB3;
  assign sine_lut64_14bit[40] = 14'h960;
  assign sine_lut64_14bit[41] = 14'h744;
  assign sine_lut64_14bit[42] = 14'h565;
  assign sine_lut64_14bit[43] = 14'h3C8;
  assign sine_lut64_14bit[44] = 14'h270;
  assign sine_lut64_14bit[45] = 14'h161;
  assign sine_lut64_14bit[46] = 14'h9E;
  assign sine_lut64_14bit[47] = 14'h28;
  assign sine_lut64_14bit[48] = 14'h1;
  assign sine_lut64_14bit[49] = 14'h28;
  assign sine_lut64_14bit[50] = 14'h9E;
  assign sine_lut64_14bit[51] = 14'h161;
  assign sine_lut64_14bit[52] = 14'h270;
  assign sine_lut64_14bit[53] = 14'h3C8;
  assign sine_lut64_14bit[54] = 14'h565;
  assign sine_lut64_14bit[55] = 14'h744;
  assign sine_lut64_14bit[56] = 14'h960;
  assign sine_lut64_14bit[57] = 14'hBB3;
  assign sine_lut64_14bit[58] = 14'hE39;
  assign sine_lut64_14bit[59] = 14'h10EA;
  assign sine_lut64_14bit[60] = 14'h13C1;
  assign sine_lut64_14bit[61] = 14'h16B6;
  assign sine_lut64_14bit[62] = 14'h19C2;
  assign sine_lut64_14bit[63] = 14'h1CDD;
